library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity fpga_project_top_level is
	generic(
		
	);
	port(
	
	);
end fpga_project_top_level;

architecture ARCH of fpga_project_top_level is

end ARCH;